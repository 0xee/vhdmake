package  c is

  constant cc : natural := 1;

end package  c;
