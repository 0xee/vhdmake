architecture b of a is

begin  -- architecture b

   
end architecture b;
