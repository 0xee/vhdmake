library ieee;
use ieee.std_logic_1164.all;

entity a is
   
  port (
    iClk : in std_ulogic);

end entity a;
